* CMOS Inverter Example for ngspice

* Power supply
VDD VDD 0 DC 5V

* Input voltage source
VIN IN 0 PWL(0 0 1n 5 2n 0 3n 5 4n 0 5n 5 6n 0)

* NMOS transistor
M1 OUT IN VSS VSS NMOS_MODEL

* PMOS transistor
M2 OUT VDD VDD VDD PMOS_MODEL

* Transistor models (simple level 1 models, replace with real models as needed)
.model NMOS_MODEL NMOS (LEVEL=1 VTO=1 KP=2.0)
.model PMOS_MODEL PMOS (LEVEL=1 VTO=-1 KP=1.0)

* Load at output (optional)
RL OUT 0 10k

* Simulation commands
.control
  run
  plot V(IN) V(OUT)
.endc

.end
