* CMOS Inverter with input and output voltage recording

* Power supplies
VDD VDD 0 DC 5V
VSS VSS 0 DC 0V

* Input voltage source (PWL waveform)
VIN IN 0 PWL(0 0 1n 5 2n 0 3n 5 4n 0 5n 5 6n 0)

* NMOS transistor
M1 OUT IN VSS VSS NMOS_MODEL

* PMOS transistor
M2 OUT VDD VDD VDD PMOS_MODEL

* Transistor models (simple level 1 models, replace with more accurate models if needed)
.model NMOS_MODEL NMOS (LEVEL=1 VTO=1 KP=2.0)
.model PMOS_MODEL PMOS (LEVEL=1 VTO=-1 KP=1.0)

* Load at output
RL OUT 0 10k

* Simulation commands
.control
  * Transient analysis for 8 ns with 10 ps timestep
  tran 10p 8n

  * Write V(IN), V(OUT), and TIME to voltages.dat
  wrdata voltages.dat V(IN) V(OUT) TIME

  quit
.endc

.end
