* CMOS Inverter with Varying Input Voltage (DC sweep)

* Power supplies
VDD VDD 0 DC 5V
VSS VSS 0 DC 0V

* Input voltage source (DC sweep)
VIN IN 0 DC 5V

* NMOS transistor
M1 OUT IN VSS VSS NMOS_MODEL

* PMOS transistor
M2 OUT VDD VDD VDD PMOS_MODEL

* Transistor models
.model NMOS_MODEL NMOS (LEVEL=1 VTO=1 KP=2.0)
.model PMOS_MODEL PMOS (LEVEL=1 VTO=-1 KP=1.0)

* Load
RL OUT 0 10k

* Simulation commands
.control
  * Sweep V(IN) from 0V to 5V in steps of 0.1V
  dc VIN 0 5 0.1

  * During the sweep, write V(IN) and V(OUT) data to voltages.dat
  wrdata voltages.dat V(IN) V(OUT)

  quit
.endc

.end
